module instruction_data_memory (
    parameter num_thirty_two_bit_words = 128;
) (
    input logic []
)